library verilog;
use verilog.vl_types.all;
entity vga_vlg_vec_tst is
end vga_vlg_vec_tst;
